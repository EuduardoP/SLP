-------------------------------------------------------------------------------
-- Title      : Porta NOT
-- Project    : Aulas de VHDL
-------------------------------------------------------------------------------
-- File       : porta_xor2.vhd
-- Author     : Giovani Baratto (gfbaratto)  <Giovani.Baratto@ufsm.br>
-- Company    : UFSM - CT - DELC
-- Created    : 2019-08-05
-- Last update: 2020-04-20
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2019-08-05  1.0      gfbaratto       Created
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
entity porta_not is
  port(x : in  std_logic;               -- entrada da porta inversora
       y : out std_logic);              -- saída da porta inversora
end entity porta_not;
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
architecture simples of porta_not is
begin
  y <= not x;
end architecture simples;
-------------------------------------------------------------------------------

