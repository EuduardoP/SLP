-------------------------------------------------------------------------------
-- Title      : Porta OR com duas entradas
-- Project    : Aulas de VHDL
-------------------------------------------------------------------------------
-- File       : porta_xor2.vhd
-- Author     : Giovani Baratto (gfbaratto)  <Giovani.Baratto@ufsm.br>
-- Company    : UFSM - CT - DELC
-- Created    : 2019-08-05
-- Last update: 2020-04-20
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2019-08-05  1.0      gfbaratto       Created
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
entity porta_or2 is
  port(x : in  std_logic;               -- uma das entradas da porta OR
       y : in  std_logic;               -- a outra entrada da porta OR
       z : out std_logic);              -- saída da porta OR
end entity porta_or2;
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
architecture simples of porta_or2 is
begin
  z <= x or y;
end architecture simples;
-------------------------------------------------------------------------------

